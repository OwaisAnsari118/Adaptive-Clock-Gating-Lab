module test();

endmodule